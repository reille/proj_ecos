# ====================================================================
#
#      i2s_stm32.cdl
#
#      eCos STM32 I2S configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      reille
# Contributors:
# Date:           2013-06-02
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_SOUND_I2S_CORTEXM_STM32 {
    display     "I2S bus driver for STM32 family of CortexM controllers"

	active_if   CYGPKG_IO
	active_if   CYGPKG_HAL_CORTEXM_STM32    
    
    include_dir cyg/io	
    description "
           This package provides a generic I2S device driver for the on-chip
           I2S peripherals in STM32 processors."

    compile     -library=libextras.a i2s_stm32.c

    define_proc {
      puts $::cdl_system_header "#define CYGDAT_DEVS_SOUND_I2S_CORTEXM_STM32_INL <cyg/io/i2s_stm32.inl>"
    }

	cdl_component CYGHWR_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2 {
		display       "ST STM32 I2S bus 2"
		active_if     { CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS2 == 0 }
		description   "
			Enable I2S bus 2 on the STM32 device.
		"
		flavor        bool
		default_value 0
		
		cdl_option CYGDAT_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2_NAME {
			display "Device name for the i2s bus2 driver for stm32"
			flavor data
			default_value {"\"/dev/i2s2\""}
			description " This option specifies the name of the i2s bus2 for stm32 
			device"
		}

		cdl_option CYGDAT_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2_MCK_ENABLE {
			display "Master clock output enable"
			flavor bool
			default_value 1
			description " This option enable master clock output"
		}

		cdl_option CYGNUM_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2_BBUF_SIZE {
			display       "Bounce buffer size"
			description   "
				DMA bounce buffers are required when running out of external
				memory.  Set this to the maximum I2S packet size which will be
				used to enable the DMA bounce buffers.  Set to 0 to disable
				bounce buffers when running from on-chip memory.
			"
			flavor        data 
			default_value 0
		}
	
		cdl_option CYGNUM_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2_DMA_TXINTR_PRI {
			display       "Transmit DMA interrupt priority"
			flavor        data
			default_value 64+7
		}

		cdl_option CYGNUM_DEVS_SOUND_I2S_CORTEXM_STM32_BUS2_DMA_RXINTR_PRI {
			display       "Receive DMA interrupt priority"
			flavor        data
			default_value 128+8
		}		
	}

	cdl_option CYGDAT_DEVS_SOUND_I2S_CORTEXM_STM32_TRACE {
		display       "Driver trace"
		flavor        bool
		default_value 0
		description   "
			Enable I2S transaction trace. Select to debug the driver."
	}
}

# EOF i2c_stm32.cdl
