# ====================================================================
#
#      mmc_stm32.cdl
#
#      MMC driver configuration data for STM32 SDIO
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      reille
# Contributors:
# Date:           2013-06-26
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_DISK_CORTEXM_STM32_MMC {
    display     "MMC driver for STM32 family of CortexM controllers"

    parent      CYGPKG_IO_DISK_DEVICES
    active_if   CYGPKG_IO_DISK
	active_if   CYGPKG_HAL_CORTEXM_STM32
    
    include_dir cyg/io	
    description "
           This package provides a MMC driver for the on-chip SDIO 
           peripherals in STM32 processors."

    compile     -library=libextras.a mmc_stm32.c


	cdl_component CYGHWR_DEVS_DISK_CORTEXM_STM32_MMC_DISK0 {
		display       "ST STM32 MMC disk 0"		
		description   "Enable the MMC disk 0 on the STM32 family of CortexM controllers."
		flavor        bool
		default_value 1
		
		cdl_option CYGDAT_DEVS_DISK_CORTEXM_STM32_MMC_DISK0_NAME {
			display "Device name for the MMC disk 0 device"
			flavor data
			default_value { "\"/dev/mmcdisk0/1\"" }
			description "
				This is the device name used to access the raw disk device
                in eCos, for example for mount operations. Note that the
                trailing slash must be present."
		}

		cdl_option CYGHWR_DEVS_DISK_CORTEXM_STM32_MMC_DISK0_DETECT_GPIO {
			display       "Card detecting GPIO"
			description   "
				This is a GPIO which are to be used to detect the card whether
				inserted or not. The GPIO is defined by the SD_DETECT_IO() 
				macro which gives the port and pin number.
			"
			flavor        data
			default_value { "SD_DETECT_IO(C, 7)" }
		}		
		
		cdl_option CYGNUM_DEVS_DISK_CORTEXM_STM32_MMC_DISK0_BBUF_SIZE {
			display       "Bounce buffer size"
			description   "
				DMA bounce buffers are required when running out of external
				memory.  Set this to the maximum SDIO packet size which will be
				used to enable the DMA bounce buffers.  Set to 0 to disable
				bounce buffers when running from on-chip memory. The value must
				be multiple of 512.
			"
			flavor        data 
			default_value 0
		}
	
		cdl_option CYGNUM_DEVS_DISK_CORTEXM_STM32_MMC_DISK0_DMA_TXINTR_PRI {
			display       "Transmit DMA interrupt priority"
			flavor        data
			default_value 64+7
		}		

		cdl_option CYGNUM_DEVS_DISK_CORTEXM_STM32_MMC_DISK0_DMA_RXINTR_PRI {
			display       "Receive DMA interrupt priority"
			flavor        data
			default_value 128+8
		}				
	}
}

# EOF mmc_stm32.cdl
