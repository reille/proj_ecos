# ====================================================================
#
#      wm8978.cdl
#
#      WM8978 - WOLFSON stereo codec with speaker driver configuration
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      reille
# Contributors:
# Date:           2013-06-02
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_SOUND_I2C_WM8978 {
    display     "WM8978 driver for WOLFSON stereo codec with speaker driver"
    
    active_if   CYGPKG_IO_FILEIO
    requires    CYGPKG_IO
    requires    CYGPKG_IO_I2C
    requires    CYGFUN_KERNEL_API_C

    include_dir cyg/io
    description "
           This package provides a sound card driver - WM8978 for 
		   WOLFSON stereo codec with speaker driver."

    define_proc {
      puts $::cdl_system_header "#define CYGDAT_DEVS_SOUND_I2C_WM8978_INL <cyg/io/wm8978.inl>"
    }
	
	compile     -library=libextras.a wm8978.c

    cdl_option CYGDAT_DEVS_SOUND_I2C_WM8978_NAME {
        display "Device name for the WM8978 driver"
        flavor data
        default_value {"\"/dev/dsp\""}
        description " This option specifies the name of the WM8978 driver 
        device"
    }

    cdl_option CYGDAT_DEVS_SOUND_I2C_WM8978_USE_I2S_DEV {
        display       "I2S channel device to used for wm8978"
        flavor        data
        default_value { "\"/dev/i2s2\"" }
        description   "
            This option selects the i2s channel device used to transact
            audio data stream with '/dev/dsp'."
    }

    cdl_option CYGDAT_DEVS_SOUND_I2C_WM8978_TRACE {
        display       "Driver trace"
        flavor        bool
        default_value 0
        description   "
            Enable wm8978 driver trace. Select to debug the driver."
    }
}

# EOF wm8978.cdl
