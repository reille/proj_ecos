# ====================================================================
#
#       stm32f10xxx_eth_driver.cdl
#
#       Ethernet driver
#       STM32F10XXX w/DM9000 platform specific support
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      reille
# Original data:  
# Contributors:   
# Date:           2013-05-10
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_CORTEXM_STM32_STM32F10XXX {
    display       "STM32F10XXX board with Davicom DM9000 ethernet driver"
    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_CORTEXM_STM32_STM32F10XXX

    include_dir   cyg/io

    # FIXME: This really belongs in the DM9000 package
    cdl_interface CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED {
        display   "Davicom DM9000 ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_DAVICOM_DM9000_INL <cyg/io/stm32f10xxx_eth_driver.inl>"
 
 	puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_DAVICOM_DM9000_CFG <pkgconf/devs_eth_cortexm_stm32_stm32f10xxx.h>"

        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }


    cdl_component CYGPKG_DEVS_ETH_CORTEXM_STM32_STM32F10XXX_ETH0 {
        display       "stm32f10xxx ethernet port driver for builtin Davicom DM9000"
        flavor        bool
        default_value 1
        description   "
            This option includes the Davicom DM9000 ethernet device driver for a
            STM32F10XXX board."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_DAVICOM_DM9000_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_CORTEXM_STM32_STM32F10XXX_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for a
                DM9000-based STM32F10XXX board."
        }
		
        cdl_option CYGDAT_DEVS_ETH_CORTEXM_STM32_STM32F10XXX_ETH0_ESA {
            display       "The ethernet station address for the ETH0 ethernet port driver"
            flavor        data
            default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
            description   "
                This option sets the ethernet station address of the ethernet device for a
                DM9000-based STM32F10XXX board."
        }		
    }



    cdl_component CYGPKG_DEVS_ETH_DM9000_ETH_REDBOOT_HOLDS_ESA {
	display         "RedBoot manages ESA initialization data"
	flavor          bool
	default_value	0

	active_if     CYGSEM_HAL_VIRTUAL_VECTOR_SUPPORT

	description   "Enabling this option will allow the ethernet
	station address to be acquired from RedBoot's configuration data,
	stored in flash memory.  It can be overridden individually by the
	'Set the ethernet station address' option for each interface."

	cdl_component CYGPKG_DEVS_ETH_DM9000_ETH_REDBOOT_HOLDS_ESA_VARS {
	    display        "Build-in flash config fields for ESAs"
	    flavor         bool
	    default_value  0

	    active_if       CYGPKG_REDBOOT
	    active_if       CYGPKG_REDBOOT_FLASH
	    active_if       CYGSEM_REDBOOT_FLASH_CONFIG
	    active_if 	    CYGPKG_REDBOOT_NETWORKING

	    description	"
	    This option controls the presence of RedBoot flash
	    configuration fields for the ESAs of the interfaces when you
	    are building RedBoot.  It is independent of whether RedBoot
	    itself uses the network or any particular interface; this
	    support is more for the application to use than for RedBoot
	    itself, though the application gets at the data by vector
	    calls; this option cannot be enabled outside of building
	    RedBoot."
	
	    cdl_option CYGVAR_ETH_DM9000_REDBOOT_HOLDS_ESA_ETH0 {
		display         "RedBoot manages ESA for eth0"
		flavor          bool
		default_value   0
	    }

            cdl_option CYGDAT_DEVS_ETH_CORTEXM_STM32_STM32F10XXX_ETH0_DEFAULT_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x00, 0x03, 0x47, 0xdf, 0x32, 0xa8}"}
                description   "The default ethernet station address. This is the
                               address used as the default value in the RedBoot
                               flash configuration field."
            }
	}
    }
}

